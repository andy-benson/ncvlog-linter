module test();
     
dda
         
         
          
    
endmodule 
