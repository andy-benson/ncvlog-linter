module lint_test();
     
dda

             
endmodule 
