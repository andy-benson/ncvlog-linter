


module test();
     
     
     woof 
     
     
     
    
endmodule 
